------- Opdracht 2/ Assignment 2 DSDL practicum
------- Altera DE10-Lite
------- ir drs E.J Boks, HAN Embedded Systems Engineering. https://ese.han.nl
------- Bibliotheek met alle componenten die in dit projekt worden gebruikt
------- Library with all components that are used in this project.

library ieee; 
use ieee.std_logic_1164.all; 

package Assignment2Package is

	component genericClockDelay is

	generic(desiredClock: integer := 10;  -- 10 Hz
           inClockFreq: natural := 100);  -- 100 Hz
			
	port 
	(
		clk,rst  : in  std_logic;
		outClock  : buffer std_logic
	);
	
	end component;
	
end Assignment2Package;
	

package body Assignment2Package is	

end Assignment2Package;



---------- 


library ieee;
use ieee.std_logic_1164.all;
use work.all;

-- Dit is een generieke klokvertraging module. Zie voorbeeld 6.2 in Pedroni 2e Editie of paragraaf 2.7 en voorbeeld 12.3 in Pedroni 3e Editie.

-- This is a generic clock delay module. See example 6.2 in Pedroni 2nd Edition or paragraph 2.7 and example 12.3 in Pedroni 3rd Edition. 

-- Maak een Test Bench aan om deze module te kunnen verifieeren.
-- Build a Test Bench in order to verify this module.
entity genericClockDelay is

	generic(desiredClock: integer := 10;  -- 10 Hz
           inClockFreq: natural := 100);  -- 100 Hz
			
	port 
	(
		clk,rst  : in  std_logic;
		outClock  : buffer std_logic
	);
	
end entity;

architecture behaviour of genericClockDelay is
	constant clockTopValue : natural := inClockFreq/(2*desiredClock);	
	
begin
	

	process (clk) 	
		variable internalCtr : natural := 0;
	begin	  
		
		if (rst ='1') then
			internalCtr := 0;
			outClock <= '0';
		elsif rising_edge(clk) then
			if internalCtr < clockTopValue then
				internalCtr := internalCtr + 1;
			else
				internalCtr := 0;
				outClock <= not outClock;
			end if;
		end if;	 
		
	end process;
	
	
end architecture;


